///////////////////////////////////////////////////////////////////////////
//                                                                       //
//			             Logarithm module [ -2.ln(x) ]                   //
//                                  By                                   //
//                        Santosh Kumar Krishnan                         //
//                                                                       //
//                         'TOP - 1' level entity                        //
//                                                                       //
///////////////////////////////////////////////////////////////////////////
/*  Copyright (C) 2016  Santosh Kumar Krishnan

    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with this program.  If not, see http://www.gnu.org/licenses/.*/
	
module log_module (
clock,
reset,
num,
value);

//input
input clock;
input reset;
input [47:0] num;

//output
output [30:0] value;

//internal registers
reg [30:0] value_d;
reg [29:0] temp_d,temp2_d;
reg [31:0] log_2_2;
reg [28:0] mul1_d;
reg [28:0] shortened_num_d1,shortened_num_dd1,shortened_num_d2,shortened_num_d3,shortened_num_d4;
reg [5:0] expo_d1,expo_d2,expo_d3,expo_d4,expo_d5,expo_d6,expo_d7;
reg [7:0] table_address_d1;
reg [18:0] c_2,c_2_d1,c_2_d2;
reg [21:0] c_1,c_1_d1,c_1_d2;
reg [29:0] c_0_t,c_0_t_d1,c_0_t_d2;
reg [18:0] ln_c_2[255:0];
reg [21:0] ln_c_1[255:0];
reg [29:0] ln_c_0[255:0];
reg [29:0] c_0_d1,c_0_d2;
reg [47:0] mul3_d; 
reg [50:0] mul2_d1,mul2_d2;
reg [37:0] expo_corr_d;
reg [33:0] adj_log_val_d;
reg [47:0] mul3_t_d;
reg [47:0] num2_d;
reg [5:0] leading_zeros_d;
reg [29:0] t1_d,t1_d1,t3_d1;
reg [28:0] t2_d;
reg [27:0] t5_d;

//internal signals
wire [47:0] num2_p1;
wire [33:0] value1;
wire [30:0] value_p;
wire [31:0] log_2_2_s;
wire [5:0] zeros_32bit;
wire [4:0] zeros_16bit;
wire [5:0] leading_zeros,leading_zeros_p1;
wire [5:0] expo,expo_p1,expo_p2,expo_p3,expo_p4,expo_p5,expo_p6,expo_p7;
wire [47:0] shifted_num;
wire [7:0] table_address,table_address_p1;
wire [18:0] c_2_p1,c_2_p2;
wire [21:0] c_1_p1,c_1_p2;
wire [29:0] c_0,c_0_p1,c_0_p2;
wire [28:0] shortened_num,shortened_num_p2,shortened_num_p1,shortened_num_pp1,shortened_num_p3,shortened_num_p4;
wire [57:0] mul1;
wire [28:0] mul1_half,mul1_half_1;
wire [50:0] mul2,mul2_p1,mul2_p2;
wire [47:0] mul3_t,mul3_t_p1;
wire [47:0] mul3,mul3_p1;
wire [29:0] temp,temp2,temp_p1,temp2_p1;
wire [30:0] log_val; 
wire log_sign;
wire [37:0] expo_corr,expo_corr_p1;
wire [33:0] adj_log_val,adj_log_val_p1; 
wire [28:0] mul1_p2;
wire [29:0] t1,t7,t8,t3,t9,t1_p1,t1_p2,t3_p1; 
wire [28:0] t2,t2_p1;
wire [27:0] t5,t6,t5_p1;
wire [29:0] c_0_t_p1,c_0_t_p2;

//combinational logic

//instantiate 16 bit leading zero detector
LZD_16 L_16_log(num[47:32],zeros_16bit);

//instantiata 32 bit leading zero detector
LZD_32 L_32_log(num[31:0],zeros_32bit);

//instantiate 48 bit left barrel shifter  
barrel_shifter_48 B_S_48(num2_p1,leading_zeros_p1,shifted_num);

//get number leading zeros and find the exponent value to be shifted by
assign leading_zeros = (zeros_16bit == 5'b10000)?(zeros_32bit + 5'b10000):zeros_16bit;

//assign values from respective flipflops.
assign num2_p1 = num2_d;
assign leading_zeros_p1 = leading_zeros_d;

//find exponent of input number.
assign expo = leading_zeros_p1 + 1;

//find address of the coefficient table
assign table_address = shifted_num[46:39];

//adjust shortened num
assign shortened_num = shifted_num[47:19];

//assign signals from respective flipflops.
assign table_address_p1 = table_address_d1;
assign shortened_num_p1 = shortened_num_d1;
assign shortened_num_pp1 = shortened_num_dd1;
assign expo_p1 = expo_d1;

//calculate the square of x in c_2*x^2-c_1*x+c_0  part 1.
assign t1 = shortened_num_pp1[28:14]*shortened_num_p1[28:14];
assign t2 = shortened_num_p1[13:0]*shortened_num_p1[28:14];
assign t5 = shortened_num_pp1[13:0]*shortened_num_pp1[13:0];

//assign signals from respective flipflops.
assign t2_p1 = t2_d;
assign t1_p1 = t1_d;
assign t5_p1 = t5_d;
assign expo_p2 = expo_d2;
assign shortened_num_p2 = shortened_num_d2;

//calculate the square of x in c_2*x^2-c_1*x+c_0  part 2.
assign t7 = {1'b0,t2_p1};
assign t6 = {15'h0,t5_p1[27:15]};
assign t8 = t7 + t6;
assign t3 = {14'b0,t8[29:13]};

//assign signals from respective flipflops.
assign t1_p2 = t1_d1;
assign t3_p1 = t3_d1;
assign shortened_num_p3 = shortened_num_d3;
assign expo_p3 = expo_d3;
assign c_0_t_p1 = c_0_t_d1;
assign c_1_p1 = c_1_d1;
assign c_2_p1 = c_2_d1;

//calculate the square of x in c_2*x^2-c_1*x+c_0  part 3.
assign t9 = t1_p2 + t3_p1;
assign mul1_half = t9[29:1];

//assign signals from respective flipflops.
assign shortened_num_p4 = shortened_num_d4;
assign mul1_p2 = mul1_d;
assign expo_p4 = expo_d4;
assign c_0_t_p2 = c_0_t_d2;
assign c_1_p2 = c_1_d2;
assign c_2_p2 = c_2_d2;

//adjust c_0
assign c_0 = {1'b0,c_0_t_p2[29:1]};

//evaluate the piecewise polynomial to find ln(shifted_num) part 1
assign mul2 = shortened_num_p4*c_1_p2;
assign mul3_t = mul1_p2*c_2_p2;

//assign signals from respective flipflops.
assign mul3_t_p1 = mul3_t_d;
assign expo_p5 = expo_d5;
assign c_0_p1 = c_0_d1;
assign mul2_p1 = mul2_d1;
 
//adjust term x*c_1 term in piecewise polynomial. 
assign mul3 = {1'b0,mul3_t_p1[47:1]};

//assign signals from respective flipflops.
assign mul3_p1 = mul3_d;
assign expo_p6 = expo_d6;
assign c_0_p2 = c_0_d2;
assign mul2_p2 = mul2_d2;

//evaluate the piecewise polynomial to find ln(shifted_num) part 2
assign temp = mul3_p1[47:18] + c_0_p2; 
assign temp2 = mul2_p2[50:21];

//assign signals from respective flipflops.
assign temp_p1 = temp_d;
assign temp2_p1 = temp2_d;
assign expo_p7 = expo_d7;

//evaluate the piecewise polynomial to find ln(shifted_num) part 3
assign log_val = temp_p1 - temp2_p1;
assign log_sign = log_val[30];

//evaluate the following ln(2)*exponent
assign log_2_2_s = log_2_2;
assign expo_corr = log_2_2_s*expo_p7;
assign adj_log_val = {log_sign,log_sign,log_sign,log_sign,log_val[29:0]};

//assign signals from respective flipflops.
assign expo_corr_p1 = expo_corr_d;
assign adj_log_val_p1 = adj_log_val_d;

//evaluate -2*ln(num) 
assign value1 = adj_log_val_p1 + expo_corr_p1[37:4]; 
assign value_p = (value1[33:31] == 3'b111)?31'h00000000:value1[33:3];

//assign value
assign value = value_d;

//sequential part

always@(posedge clock)
begin
//reset = 0? update all the registers.
	if(reset == 1'b0)
	begin
		log_2_2 = 32'hB17217F7;
		value_d = value_p;
		expo_corr_d = expo_corr;
		leading_zeros_d = leading_zeros;
		num2_d = num;
		expo_d1 = expo;
		expo_d2 = expo_p1;
		expo_d3 = expo_p2;
		expo_d4 = expo_p3;
		expo_d5 = expo_p4;
		expo_d6 = expo_p5;
		expo_d7 = expo_p6;
		t1_d = t1;
		t2_d = t2;
		t5_d = t5;
		t3_d1 = t3;
		t1_d1 = t1_p1;
		c_0_t_d1 = c_0_t;
		c_1_d1 = c_1;
		c_2_d1 = c_2;
		c_0_t_d2 = c_0_t_p1;
        c_1_d2 = c_1_p1;
        c_2_d2 = c_2_p1;
		temp_d = temp;
		temp2_d = temp2;
		c_0_d1 = c_0;
		c_0_d2 = c_0_p1;
		mul2_d1 = mul2;
		mul2_d2 = mul2_p1;
		mul3_d = mul3;
	    mul3_t_d = mul3_t;
		adj_log_val_d = adj_log_val;
		shortened_num_d1 = shortened_num;
		shortened_num_dd1 = shortened_num;
		shortened_num_d2 = shortened_num_p1;
		shortened_num_d3 = shortened_num_p2;
		shortened_num_d4 = shortened_num_p3;
		table_address_d1 = table_address;
		mul1_d = mul1_half;
		ln_c_2[0] = 19'h7F807;
		ln_c_2[1] = 19'h7E836;
		ln_c_2[2] = 19'h7D895;
		ln_c_2[3] = 19'h7C921;
		ln_c_2[4] = 19'h7B9DC;
		ln_c_2[5] = 19'h7AAC2;
		ln_c_2[6] = 19'h79BD5;
		ln_c_2[7] = 19'h78D14;
		ln_c_2[8] = 19'h77E7D;
		ln_c_2[9] = 19'h77010;
		ln_c_2[10] = 19'h761CD;
		ln_c_2[11] = 19'h753B3;
		ln_c_2[12] = 19'h745C0;
		ln_c_2[13] = 19'h737F6;
		ln_c_2[14] = 19'h72A53;
		ln_c_2[15] = 19'h71CD6;
		ln_c_2[16] = 19'h70F7F;
		ln_c_2[17] = 19'h7024D;
		ln_c_2[18] = 19'h6F541;
		ln_c_2[19] = 19'h6E858;
		ln_c_2[20] = 19'h6DB94;
		ln_c_2[21] = 19'h6CEF3;
		ln_c_2[22] = 19'h6C274;
		ln_c_2[23] = 19'h6B618;
		ln_c_2[24] = 19'h6A9DD;
		ln_c_2[25] = 19'h69DC4;
		ln_c_2[26] = 19'h691CC;
		ln_c_2[27] = 19'h685F4;
		ln_c_2[28] = 19'h67A3C;
		ln_c_2[29] = 19'h66EA3;
		ln_c_2[30] = 19'h6632A;
		ln_c_2[31] = 19'h657CF;
		ln_c_2[32] = 19'h64C92;
		ln_c_2[33] = 19'h64173;
		ln_c_2[34] = 19'h63671;
		ln_c_2[35] = 19'h62B8C;
		ln_c_2[36] = 19'h620C4;
		ln_c_2[37] = 19'h61618;
		ln_c_2[38] = 19'h60B88;
		ln_c_2[39] = 19'h60113;
		ln_c_2[40] = 19'h5F6B9;
		ln_c_2[41] = 19'h5EC7A;
		ln_c_2[42] = 19'h5E256;
		ln_c_2[43] = 19'h5D84B;
		ln_c_2[44] = 19'h5CE5A;
		ln_c_2[45] = 19'h5C482;
		ln_c_2[46] = 19'h5BAC3;
		ln_c_2[47] = 19'h5B11C;
		ln_c_2[48] = 19'h5A78E;
		ln_c_2[49] = 19'h59E18;
		ln_c_2[50] = 19'h594BA;
		ln_c_2[51] = 19'h58B73;
		ln_c_2[52] = 19'h58243;
		ln_c_2[53] = 19'h5792A;
		ln_c_2[54] = 19'h57027;
		ln_c_2[55] = 19'h5673A;
		ln_c_2[56] = 19'h55E64;
		ln_c_2[57] = 19'h555A3;
		ln_c_2[58] = 19'h54CF7;
		ln_c_2[59] = 19'h54460;
		ln_c_2[60] = 19'h53BDF;
		ln_c_2[61] = 19'h53371;
		ln_c_2[62] = 19'h52B18;
		ln_c_2[63] = 19'h522D3;
		ln_c_2[64] = 19'h51AA2;
		ln_c_2[65] = 19'h51285;
		ln_c_2[66] = 19'h50A7A;
		ln_c_2[67] = 19'h50283;
		ln_c_2[68] = 19'h4FA9F;
		ln_c_2[69] = 19'h4F2CD;
		ln_c_2[70] = 19'h4EB0D;
		ln_c_2[71] = 19'h4E360;
		ln_c_2[72] = 19'h4DBC4;
		ln_c_2[73] = 19'h4D43B;
		ln_c_2[74] = 19'h4CCC2;
		ln_c_2[75] = 19'h4C55B;
		ln_c_2[76] = 19'h4BE06;
		ln_c_2[77] = 19'h4B6C1;
		ln_c_2[78] = 19'h4AF8C;
		ln_c_2[79] = 19'h4A868;
		ln_c_2[80] = 19'h4A155;
		ln_c_2[81] = 19'h49A51;
		ln_c_2[82] = 19'h4935E;
		ln_c_2[83] = 19'h48C7A;
		ln_c_2[84] = 19'h485A5;
		ln_c_2[85] = 19'h47EE0;
		ln_c_2[86] = 19'h4782A;
		ln_c_2[87] = 19'h47183;
		ln_c_2[88] = 19'h46AEB;
		ln_c_2[89] = 19'h46462;
		ln_c_2[90] = 19'h45DE7;
		ln_c_2[91] = 19'h4577A;
		ln_c_2[92] = 19'h4511B;
		ln_c_2[93] = 19'h44ACB;
		ln_c_2[94] = 19'h44488;
		ln_c_2[95] = 19'h43E53;
		ln_c_2[96] = 19'h4382B;
		ln_c_2[97] = 19'h43211;
		ln_c_2[98] = 19'h42C04;
		ln_c_2[99] = 19'h42604;
		ln_c_2[100] = 19'h42011;
		ln_c_2[101] = 19'h41A2A;
		ln_c_2[102] = 19'h41450;
		ln_c_2[103] = 19'h40E83;
		ln_c_2[104] = 19'h408C2;
		ln_c_2[105] = 19'h4030E;
		ln_c_2[106] = 19'h3FD65;
		ln_c_2[107] = 19'h3F7C8;
		ln_c_2[108] = 19'h3F237;
		ln_c_2[109] = 19'h3ECB2;
		ln_c_2[110] = 19'h3E739;
		ln_c_2[111] = 19'h3E1CA;
		ln_c_2[112] = 19'h3DC67;
		ln_c_2[113] = 19'h3D710;
		ln_c_2[114] = 19'h3D1C3;
		ln_c_2[115] = 19'h3CC81;
		ln_c_2[116] = 19'h3C74A;
		ln_c_2[117] = 19'h3C21E;
		ln_c_2[118] = 19'h3BCFD;
		ln_c_2[119] = 19'h3B7E5;
		ln_c_2[120] = 19'h3B2D9;
		ln_c_2[121] = 19'h3ADD6;
		ln_c_2[122] = 19'h3A8DE;
		ln_c_2[123] = 19'h3A3F0;
		ln_c_2[124] = 19'h39F0B;
		ln_c_2[125] = 19'h39A31;
		ln_c_2[126] = 19'h39560;
		ln_c_2[127] = 19'h39099;
		ln_c_2[128] = 19'h38BDB;
		ln_c_2[129] = 19'h38727;
		ln_c_2[130] = 19'h3827C;
		ln_c_2[131] = 19'h37DDA;
		ln_c_2[132] = 19'h37942;
		ln_c_2[133] = 19'h374B2;
		ln_c_2[134] = 19'h3702C;
		ln_c_2[135] = 19'h36BAE;
		ln_c_2[136] = 19'h36739;
		ln_c_2[137] = 19'h362CD;
		ln_c_2[138] = 19'h35E6A;
		ln_c_2[139] = 19'h35A0F;
		ln_c_2[140] = 19'h355BC;
		ln_c_2[141] = 19'h35172;
		ln_c_2[142] = 19'h34D30;
		ln_c_2[143] = 19'h348F6;
		ln_c_2[144] = 19'h344C4;
		ln_c_2[145] = 19'h3409A;
		ln_c_2[146] = 19'h33C79;
		ln_c_2[147] = 19'h3385F;
		ln_c_2[148] = 19'h3344D;
		ln_c_2[149] = 19'h33042;
		ln_c_2[150] = 19'h32C3F;
		ln_c_2[151] = 19'h32844;
		ln_c_2[152] = 19'h32450;
		ln_c_2[153] = 19'h32064;
		ln_c_2[154] = 19'h31C7F;
		ln_c_2[155] = 19'h318A1;
		ln_c_2[156] = 19'h314CA;
		ln_c_2[157] = 19'h310FB;
		ln_c_2[158] = 19'h30D32;
		ln_c_2[159] = 19'h30971;
		ln_c_2[160] = 19'h305B6;
		ln_c_2[161] = 19'h30202;
		ln_c_2[162] = 19'h2FE56;
		ln_c_2[163] = 19'h2FAAF;
		ln_c_2[164] = 19'h2F710;
		ln_c_2[165] = 19'h2F377;
		ln_c_2[166] = 19'h2EFE4;
		ln_c_2[167] = 19'h2EC59;
		ln_c_2[168] = 19'h2E8D3;
		ln_c_2[169] = 19'h2E554;
		ln_c_2[170] = 19'h2E1DB;
		ln_c_2[171] = 19'h2DE68;
		ln_c_2[172] = 19'h2DAFC;
		ln_c_2[173] = 19'h2D795;
		ln_c_2[174] = 19'h2D435;
		ln_c_2[175] = 19'h2D0DB;
		ln_c_2[176] = 19'h2CD86;
		ln_c_2[177] = 19'h2CA38;
		ln_c_2[178] = 19'h2C6EF;
		ln_c_2[179] = 19'h2C3AC;
		ln_c_2[180] = 19'h2C06F;
		ln_c_2[181] = 19'h2BD38;
		ln_c_2[182] = 19'h2BA06;
		ln_c_2[183] = 19'h2B6DA;
		ln_c_2[184] = 19'h2B3B3;
		ln_c_2[185] = 19'h2B092;
		ln_c_2[186] = 19'h2AD76;
		ln_c_2[187] = 19'h2AA5F;
		ln_c_2[188] = 19'h2A74E;
		ln_c_2[189] = 19'h2A443;
		ln_c_2[190] = 19'h2A13C;
		ln_c_2[191] = 19'h29E3A;
		ln_c_2[192] = 19'h29B3E;
		ln_c_2[193] = 19'h29847;
		ln_c_2[194] = 19'h29555;
		ln_c_2[195] = 19'h29268;
		ln_c_2[196] = 19'h28F80;
		ln_c_2[197] = 19'h28C9C;
		ln_c_2[198] = 19'h289BE;
		ln_c_2[199] = 19'h286E4;
		ln_c_2[200] = 19'h28410;
		ln_c_2[201] = 19'h28140;
		ln_c_2[202] = 19'h27E74;
		ln_c_2[203] = 19'h27BAE;
		ln_c_2[204] = 19'h278EC;
		ln_c_2[205] = 19'h2762E;
		ln_c_2[206] = 19'h27376;
		ln_c_2[207] = 19'h270C1;
		ln_c_2[208] = 19'h26E11;
		ln_c_2[209] = 19'h26B66;
		ln_c_2[210] = 19'h268BF;
		ln_c_2[211] = 19'h2661C;
		ln_c_2[212] = 19'h2637E;
		ln_c_2[213] = 19'h260E3;
		ln_c_2[214] = 19'h25E4E;
		ln_c_2[215] = 19'h25BBC;
		ln_c_2[216] = 19'h2592E;
		ln_c_2[217] = 19'h256A5;
		ln_c_2[218] = 19'h25420;
		ln_c_2[219] = 19'h2519E;
		ln_c_2[220] = 19'h24F21;
		ln_c_2[221] = 19'h24CA8;
		ln_c_2[222] = 19'h24A33;
		ln_c_2[223] = 19'h247C2;
		ln_c_2[224] = 19'h24554;
		ln_c_2[225] = 19'h242EB;
		ln_c_2[226] = 19'h24085;
		ln_c_2[227] = 19'h23E23;
		ln_c_2[228] = 19'h23BC5;
		ln_c_2[229] = 19'h2396B;
		ln_c_2[230] = 19'h23714;
		ln_c_2[231] = 19'h234C1;
		ln_c_2[232] = 19'h23272;
		ln_c_2[233] = 19'h23026;
		ln_c_2[234] = 19'h22DDE;
		ln_c_2[235] = 19'h22B99;
		ln_c_2[236] = 19'h22958;
		ln_c_2[237] = 19'h2271B;
		ln_c_2[238] = 19'h224E1;
		ln_c_2[239] = 19'h222AA;
		ln_c_2[240] = 19'h22077;
		ln_c_2[241] = 19'h21E47;
		ln_c_2[242] = 19'h21C1B;
		ln_c_2[243] = 19'h219F2;
		ln_c_2[244] = 19'h217CC;
		ln_c_2[245] = 19'h215AA;
		ln_c_2[246] = 19'h2138A;
		ln_c_2[247] = 19'h2116E;
		ln_c_2[248] = 19'h20F56;
		ln_c_2[249] = 19'h20D40;
		ln_c_2[250] = 19'h20B2E;
		ln_c_2[251] = 19'h2091E;
		ln_c_2[252] = 19'h20712;
		ln_c_2[253] = 19'h20509;
		ln_c_2[254] = 19'h20303;
		ln_c_2[255] = 19'h20100;

		ln_c_1[0] = 22'h3FE016;
		ln_c_1[1] = 22'h3FA096;
		ln_c_1[2] = 22'h3F6192;
		ln_c_1[3] = 22'h3F230C;
		ln_c_1[4] = 22'h3EE500;
		ln_c_1[5] = 22'h3EA76D;
		ln_c_1[6] = 22'h3E6A53;
		ln_c_1[7] = 22'h3E2DAF;
		ln_c_1[8] = 22'h3DF181;
		ln_c_1[9] = 22'h3DB5C7;
		ln_c_1[10] = 22'h3D7A80;
		ln_c_1[11] = 22'h3D3FAA;
		ln_c_1[12] = 22'h3D0544;
		ln_c_1[13] = 22'h3CCB4D;
		ln_c_1[14] = 22'h3C91C4;
		ln_c_1[15] = 22'h3C58A8;
		ln_c_1[16] = 22'h3C1FF6;
		ln_c_1[17] = 22'h3BE7AF;
		ln_c_1[18] = 22'h3BAFD1;
		ln_c_1[19] = 22'h3B785B;
		ln_c_1[20] = 22'h3B414B;
		ln_c_1[21] = 22'h3B0AA1;
		ln_c_1[22] = 22'h3AD45B;
		ln_c_1[23] = 22'h3A9E79;
		ln_c_1[24] = 22'h3A68F9;
		ln_c_1[25] = 22'h3A33DB;
		ln_c_1[26] = 22'h39FF1D;
		ln_c_1[27] = 22'h39CABE;
		ln_c_1[28] = 22'h3996BD;
		ln_c_1[29] = 22'h39631A;
		ln_c_1[30] = 22'h392FD2;
		ln_c_1[31] = 22'h38FCE7;
		ln_c_1[32] = 22'h38CA55;
		ln_c_1[33] = 22'h38981D;
		ln_c_1[34] = 22'h38663E;
		ln_c_1[35] = 22'h3834B6;
		ln_c_1[36] = 22'h380384;
		ln_c_1[37] = 22'h37D2A9;
		ln_c_1[38] = 22'h37A223;
		ln_c_1[39] = 22'h3771F0;
		ln_c_1[40] = 22'h374211;
		ln_c_1[41] = 22'h371284;
		ln_c_1[42] = 22'h36E349;
		ln_c_1[43] = 22'h36B45E;
		ln_c_1[44] = 22'h3685C4;
		ln_c_1[45] = 22'h365779;
		ln_c_1[46] = 22'h36297B;
		ln_c_1[47] = 22'h35FBCC;
		ln_c_1[48] = 22'h35CE69;
		ln_c_1[49] = 22'h35A153;
		ln_c_1[50] = 22'h357488;
		ln_c_1[51] = 22'h354807;
		ln_c_1[52] = 22'h351BD0;
		ln_c_1[53] = 22'h34EFE2;
		ln_c_1[54] = 22'h34C43D;
		ln_c_1[55] = 22'h3498E0;
		ln_c_1[56] = 22'h346DC9;
		ln_c_1[57] = 22'h3442F9;
		ln_c_1[58] = 22'h34186F;
		ln_c_1[59] = 22'h33EE29;
		ln_c_1[60] = 22'h33C428;
		ln_c_1[61] = 22'h339A6B;
		ln_c_1[62] = 22'h3370F1;
		ln_c_1[63] = 22'h3347B9;
		ln_c_1[64] = 22'h331EC4;
		ln_c_1[65] = 22'h32F60F;
		ln_c_1[66] = 22'h32CD9B;
		ln_c_1[67] = 22'h32A567;
		ln_c_1[68] = 22'h327D73;
		ln_c_1[69] = 22'h3255BD;
		ln_c_1[70] = 22'h322E46;
		ln_c_1[71] = 22'h32070C;
		ln_c_1[72] = 22'h31E00F;
		ln_c_1[73] = 22'h31B94F;
		ln_c_1[74] = 22'h3192CB;
		ln_c_1[75] = 22'h316C83;
		ln_c_1[76] = 22'h314675;
		ln_c_1[77] = 22'h3120A2;
		ln_c_1[78] = 22'h30FB09;
		ln_c_1[79] = 22'h30D5A9;
		ln_c_1[80] = 22'h30B082;
		ln_c_1[81] = 22'h308B94;
		ln_c_1[82] = 22'h3066DD;
		ln_c_1[83] = 22'h30425E;
		ln_c_1[84] = 22'h301E15;
		ln_c_1[85] = 22'h2FFA03;
		ln_c_1[86] = 22'h2FD627;
		ln_c_1[87] = 22'h2FB280;
		ln_c_1[88] = 22'h2F8F0F;
		ln_c_1[89] = 22'h2F6BD1;
		ln_c_1[90] = 22'h2F48C8;
		ln_c_1[91] = 22'h2F25F3;
		ln_c_1[92] = 22'h2F0351;
		ln_c_1[93] = 22'h2EE0E1;
		ln_c_1[94] = 22'h2EBEA4;
		ln_c_1[95] = 22'h2E9C98;
		ln_c_1[96] = 22'h2E7ABE;
		ln_c_1[97] = 22'h2E5915;
		ln_c_1[98] = 22'h2E379D;
		ln_c_1[99] = 22'h2E1655;
		ln_c_1[100] = 22'h2DF53D;
		ln_c_1[101] = 22'h2DD454;
		ln_c_1[102] = 22'h2DB39A;
		ln_c_1[103] = 22'h2D930E;
		ln_c_1[104] = 22'h2D72B1;
		ln_c_1[105] = 22'h2D5282;
		ln_c_1[106] = 22'h2D3280;
		ln_c_1[107] = 22'h2D12AC;
		ln_c_1[108] = 22'h2CF304;
		ln_c_1[109] = 22'h2CD388;
		ln_c_1[110] = 22'h2CB438;
		ln_c_1[111] = 22'h2C9514;
		ln_c_1[112] = 22'h2C761C;
		ln_c_1[113] = 22'h2C574E;
		ln_c_1[114] = 22'h2C38AA;
		ln_c_1[115] = 22'h2C1A31;
		ln_c_1[116] = 22'h2BFBE2;
		ln_c_1[117] = 22'h2BDDBD;
		ln_c_1[118] = 22'h2BBFC0;
		ln_c_1[119] = 22'h2BA1ED;
		ln_c_1[120] = 22'h2B8442;
		ln_c_1[121] = 22'h2B66BF;
		ln_c_1[122] = 22'h2B4964;
		ln_c_1[123] = 22'h2B2C31;
		ln_c_1[124] = 22'h2B0F25;
		ln_c_1[125] = 22'h2AF240;
		ln_c_1[126] = 22'h2AD582;
		ln_c_1[127] = 22'h2AB8EA;
		ln_c_1[128] = 22'h2A9C78;
		ln_c_1[129] = 22'h2A802C;
		ln_c_1[130] = 22'h2A6406;
		ln_c_1[131] = 22'h2A4804;
		ln_c_1[132] = 22'h2A2C28;
		ln_c_1[133] = 22'h2A1070;
		ln_c_1[134] = 22'h29F4DC;
		ln_c_1[135] = 22'h29D96D;
		ln_c_1[136] = 22'h29BE21;
		ln_c_1[137] = 22'h29A2F9;
		ln_c_1[138] = 22'h2987F4;
		ln_c_1[139] = 22'h296D13;
		ln_c_1[140] = 22'h295253;
		ln_c_1[141] = 22'h2937B7;
		ln_c_1[142] = 22'h291D3C;
		ln_c_1[143] = 22'h2902E4;
		ln_c_1[144] = 22'h28E8AD;
		ln_c_1[145] = 22'h28CE97;
		ln_c_1[146] = 22'h28B4A3;
		ln_c_1[147] = 22'h289ACF;
		ln_c_1[148] = 22'h28811D;
		ln_c_1[149] = 22'h28678B;
		ln_c_1[150] = 22'h284E19;
		ln_c_1[151] = 22'h2834C6;
		ln_c_1[152] = 22'h281B94;
		ln_c_1[153] = 22'h280281;
		ln_c_1[154] = 22'h27E98E;
		ln_c_1[155] = 22'h27D0B9;
		ln_c_1[156] = 22'h27B804;
		ln_c_1[157] = 22'h279F6D;
		ln_c_1[158] = 22'h2786F4;
		ln_c_1[159] = 22'h276E99;
		ln_c_1[160] = 22'h27565D;
		ln_c_1[161] = 22'h273E3E;
		ln_c_1[162] = 22'h27263C;
		ln_c_1[163] = 22'h270E58;
		ln_c_1[164] = 22'h26F691;
		ln_c_1[165] = 22'h26DEE7;
		ln_c_1[166] = 22'h26C75A;
		ln_c_1[167] = 22'h26AFE9;
		ln_c_1[168] = 22'h269894;
		ln_c_1[169] = 22'h26815C;
		ln_c_1[170] = 22'h266A3F;
		ln_c_1[171] = 22'h26533E;
		ln_c_1[172] = 22'h263C58;
		ln_c_1[173] = 22'h26258E;
		ln_c_1[174] = 22'h260EDF;
		ln_c_1[175] = 22'h25F84B;
		ln_c_1[176] = 22'h25E1D1;
		ln_c_1[177] = 22'h25CB72;
		ln_c_1[178] = 22'h25B52D;
		ln_c_1[179] = 22'h259F03;
		ln_c_1[180] = 22'h2588F3;
		ln_c_1[181] = 22'h2572FC;
		ln_c_1[182] = 22'h255D1F;
		ln_c_1[183] = 22'h25475B;
		ln_c_1[184] = 22'h2531B1;
		ln_c_1[185] = 22'h251C20;
		ln_c_1[186] = 22'h2506A8;
		ln_c_1[187] = 22'h24F149;
		ln_c_1[188] = 22'h24DC02;
		ln_c_1[189] = 22'h24C6D4;
		ln_c_1[190] = 22'h24B1BE;
		ln_c_1[191] = 22'h249CC0;
		ln_c_1[192] = 22'h2487DA;
		ln_c_1[193] = 22'h24730C;
		ln_c_1[194] = 22'h245E55;
		ln_c_1[195] = 22'h2449B6;
		ln_c_1[196] = 22'h24352F;
		ln_c_1[197] = 22'h2420BE;
		ln_c_1[198] = 22'h240C65;
		ln_c_1[199] = 22'h23F822;
		ln_c_1[200] = 22'h23E3F7;
		ln_c_1[201] = 22'h23CFE1;
		ln_c_1[202] = 22'h23BBE3;
		ln_c_1[203] = 22'h23A7FA;
		ln_c_1[204] = 22'h239428;
		ln_c_1[205] = 22'h23806B;
		ln_c_1[206] = 22'h236CC5;
		ln_c_1[207] = 22'h235934;
		ln_c_1[208] = 22'h2345B8;
		ln_c_1[209] = 22'h233253;
		ln_c_1[210] = 22'h231F02;
		ln_c_1[211] = 22'h230BC7;
		ln_c_1[212] = 22'h22F8A0;
		ln_c_1[213] = 22'h22E58F;
		ln_c_1[214] = 22'h22D292;
		ln_c_1[215] = 22'h22BFAA;
		ln_c_1[216] = 22'h22ACD6;
		ln_c_1[217] = 22'h229A17;
		ln_c_1[218] = 22'h22876C;
		ln_c_1[219] = 22'h2274D5;
		ln_c_1[220] = 22'h226252;
		ln_c_1[221] = 22'h224FE3;
		ln_c_1[222] = 22'h223D87;
		ln_c_1[223] = 22'h222B3F;
		ln_c_1[224] = 22'h22190B;
		ln_c_1[225] = 22'h2206EA;
		ln_c_1[226] = 22'h21F4DC;
		ln_c_1[227] = 22'h21E2E2;
		ln_c_1[228] = 22'h21D0FA;
		ln_c_1[229] = 22'h21BF25;
		ln_c_1[230] = 22'h21AD63;
		ln_c_1[231] = 22'h219BB4;
		ln_c_1[232] = 22'h218A17;
		ln_c_1[233] = 22'h21788D;
		ln_c_1[234] = 22'h216715;
		ln_c_1[235] = 22'h2155AF;
		ln_c_1[236] = 22'h21445B;
		ln_c_1[237] = 22'h213319;
		ln_c_1[238] = 22'h2121E9;
		ln_c_1[239] = 22'h2110CB;
		ln_c_1[240] = 22'h20FFBE;
		ln_c_1[241] = 22'h20EEC3;
		ln_c_1[242] = 22'h20DDDA;
		ln_c_1[243] = 22'h20CD02;
		ln_c_1[244] = 22'h20BC3B;
		ln_c_1[245] = 22'h20AB85;
		ln_c_1[246] = 22'h209AE0;
		ln_c_1[247] = 22'h208A4C;
		ln_c_1[248] = 22'h2079C9;
		ln_c_1[249] = 22'h206957;
		ln_c_1[250] = 22'h2058F5;
		ln_c_1[251] = 22'h2048A4;
		ln_c_1[252] = 22'h203863;
		ln_c_1[253] = 22'h202833;
		ln_c_1[254] = 22'h201812;
		ln_c_1[255] = 22'h200802;

		ln_c_0[0] = 30'h2FF0087A;
		ln_c_0[1] = 30'h2FD0284F;
		ln_c_0[2] = 30'h2FB067C3;
		ln_c_0[3] = 30'h2F90C69B;
		ln_c_0[4] = 30'h2F714498;
		ln_c_0[5] = 30'h2F51E17D;
		ln_c_0[6] = 30'h2F329D0C;
		ln_c_0[7] = 30'h2F13770B;
		ln_c_0[8] = 30'h2EF46F3F;
		ln_c_0[9] = 30'h2ED5856C;
		ln_c_0[10] = 30'h2EB6B95B;
		ln_c_0[11] = 30'h2E980ACF;
		ln_c_0[12] = 30'h2E797994;
		ln_c_0[13] = 30'h2E5B056F;
		ln_c_0[14] = 30'h2E3CAE2B;
		ln_c_0[15] = 30'h2E1E738E;
		ln_c_0[16] = 30'h2E005567;
		ln_c_0[17] = 30'h2DE2537D;
		ln_c_0[18] = 30'h2DC46D9D;
		ln_c_0[19] = 30'h2DA6A391;
		ln_c_0[20] = 30'h2D88F528;
		ln_c_0[21] = 30'h2D6B622C;
		ln_c_0[22] = 30'h2D4DEA6D;
		ln_c_0[23] = 30'h2D308DB8;
		ln_c_0[24] = 30'h2D134BDA;
		ln_c_0[25] = 30'h2CF624A5;
		ln_c_0[26] = 30'h2CD917E7;
		ln_c_0[27] = 30'h2CBC2570;
		ln_c_0[28] = 30'h2C9F4D10;
		ln_c_0[29] = 30'h2C828E9B;
		ln_c_0[30] = 30'h2C65E9DF;
		ln_c_0[31] = 30'h2C495EB1;
		ln_c_0[32] = 30'h2C2CECE2;
		ln_c_0[33] = 30'h2C109444;
		ln_c_0[34] = 30'h2BF454AD;
		ln_c_0[35] = 30'h2BD82DF0;
		ln_c_0[36] = 30'h2BBC1FE1;
		ln_c_0[37] = 30'h2BA02A56;
		ln_c_0[38] = 30'h2B844D23;
		ln_c_0[39] = 30'h2B68881E;
		ln_c_0[40] = 30'h2B4CDB1D;
		ln_c_0[41] = 30'h2B3145F8;
		ln_c_0[42] = 30'h2B15C883;
		ln_c_0[43] = 30'h2AFA6299;
		ln_c_0[44] = 30'h2ADF1410;
		ln_c_0[45] = 30'h2AC3DCC1;
		ln_c_0[46] = 30'h2AA8BC84;
		ln_c_0[47] = 30'h2A8DB331;
		ln_c_0[48] = 30'h2A72C0A4;
		ln_c_0[49] = 30'h2A57E4B4;
		ln_c_0[50] = 30'h2A3D1F3D;
		ln_c_0[51] = 30'h2A22701A;
		ln_c_0[52] = 30'h2A07D723;
		ln_c_0[53] = 30'h29ED5436;
		ln_c_0[54] = 30'h29D2E72E;
		ln_c_0[55] = 30'h29B88FE6;
		ln_c_0[56] = 30'h299E4E3B;
		ln_c_0[57] = 30'h2984220C;
		ln_c_0[58] = 30'h296A0B31;
		ln_c_0[59] = 30'h2950098A;
		ln_c_0[60] = 30'h29361CF5;
		ln_c_0[61] = 30'h291C4550;
		ln_c_0[62] = 30'h29028278;
		ln_c_0[63] = 30'h28E8D44E;
		ln_c_0[64] = 30'h28CF3AAF;
		ln_c_0[65] = 30'h28B5B57A;
		ln_c_0[66] = 30'h289C448E;
		ln_c_0[67] = 30'h2882E7CD;
		ln_c_0[68] = 30'h28699F17;
		ln_c_0[69] = 30'h28506A4B;
		ln_c_0[70] = 30'h2837494A;
		ln_c_0[71] = 30'h281E3BF6;
		ln_c_0[72] = 30'h2805422D;
		ln_c_0[73] = 30'h27EC5BD7;
		ln_c_0[74] = 30'h27D388CF;
		ln_c_0[75] = 30'h27BAC8FC;
		ln_c_0[76] = 30'h27A21C3D;
		ln_c_0[77] = 30'h27898277;
		ln_c_0[78] = 30'h2770FB8B;
		ln_c_0[79] = 30'h2758875E;
		ln_c_0[80] = 30'h274025D2;
		ln_c_0[81] = 30'h2727D6CE;
		ln_c_0[82] = 30'h270F9A31;
		ln_c_0[83] = 30'h26F76FE1;
		ln_c_0[84] = 30'h26DF57C5;
		ln_c_0[85] = 30'h26C751BE;
		ln_c_0[86] = 30'h26AF5DB3;
		ln_c_0[87] = 30'h26977B8A;
		ln_c_0[88] = 30'h267FAB25;
		ln_c_0[89] = 30'h2667EC6C;
		ln_c_0[90] = 30'h26503F45;
		ln_c_0[91] = 30'h2638A397;
		ln_c_0[92] = 30'h26211946;
		ln_c_0[93] = 30'h2609A039;
		ln_c_0[94] = 30'h25F23858;
		ln_c_0[95] = 30'h25DAE189;
		ln_c_0[96] = 30'h25C39BB3;
		ln_c_0[97] = 30'h25AC66BD;
		ln_c_0[98] = 30'h25954290;
		ln_c_0[99] = 30'h257E2F13;
		ln_c_0[100] = 30'h25672C2E;
		ln_c_0[101] = 30'h255039CA;
		ln_c_0[102] = 30'h253957CF;
		ln_c_0[103] = 30'h25228625;
		ln_c_0[104] = 30'h250BC4B5;
		ln_c_0[105] = 30'h24F51367;
		ln_c_0[106] = 30'h24DE7225;
		ln_c_0[107] = 30'h24C7E0DA;
		ln_c_0[108] = 30'h24B15F6E;
		ln_c_0[109] = 30'h249AEDCB;
		ln_c_0[110] = 30'h24848BDB;
		ln_c_0[111] = 30'h246E3987;
		ln_c_0[112] = 30'h2457F6BC;
		ln_c_0[113] = 30'h2441C360;
		ln_c_0[114] = 30'h242B9F63;
		ln_c_0[115] = 30'h24158AAB;
		ln_c_0[116] = 30'h23FF8526;
		ln_c_0[117] = 30'h23E98EBE;
		ln_c_0[118] = 30'h23D3A75E;
		ln_c_0[119] = 30'h23BDCEF3;
		ln_c_0[120] = 30'h23A80567;
		ln_c_0[121] = 30'h23924AA6;
		ln_c_0[122] = 30'h237C9E9D;
		ln_c_0[123] = 30'h23670138;
		ln_c_0[124] = 30'h23517263;
		ln_c_0[125] = 30'h233BF209;
		ln_c_0[126] = 30'h23268017;
		ln_c_0[127] = 30'h23111C7D;
		ln_c_0[128] = 30'h22FBC724;
		ln_c_0[129] = 30'h22E67FFB;
		ln_c_0[130] = 30'h22D146EF;
		ln_c_0[131] = 30'h22BC1BEB;
		ln_c_0[132] = 30'h22A6FEE0;
		ln_c_0[133] = 30'h2291EFB9;
		ln_c_0[134] = 30'h227CEE67;
		ln_c_0[135] = 30'h2267FAD4;
		ln_c_0[136] = 30'h225314EF;
		ln_c_0[137] = 30'h223E3CA8;
		ln_c_0[138] = 30'h222971ED;
		ln_c_0[139] = 30'h2214B4AA;
		ln_c_0[140] = 30'h220004D1;
		ln_c_0[141] = 30'h21EB624E;
		ln_c_0[142] = 30'h21D6CD12;
		ln_c_0[143] = 30'h21C24509;
		ln_c_0[144] = 30'h21ADCA24;
		ln_c_0[145] = 30'h21995C53;
		ln_c_0[146] = 30'h2184FB85;
		ln_c_0[147] = 30'h2170A7A7;
		ln_c_0[148] = 30'h215C60AD;
		ln_c_0[149] = 30'h21482683;
		ln_c_0[150] = 30'h2133F91A;
		ln_c_0[151] = 30'h211FD862;
		ln_c_0[152] = 30'h210BC44A;
		ln_c_0[153] = 30'h20F7BCC5;
		ln_c_0[154] = 30'h20E3C1C0;
		ln_c_0[155] = 30'h20CFD32E;
		ln_c_0[156] = 30'h20BBF0FF;
		ln_c_0[157] = 30'h20A81B22;
		ln_c_0[158] = 30'h2094518B;
		ln_c_0[159] = 30'h20809426;
		ln_c_0[160] = 30'h206CE2E9;
		ln_c_0[161] = 30'h20593DC2;
		ln_c_0[162] = 30'h2045A4A3;
		ln_c_0[163] = 30'h2032177E;
		ln_c_0[164] = 30'h201E9643;
		ln_c_0[165] = 30'h200B20E4;
		ln_c_0[166] = 30'h1FF7B755;
		ln_c_0[167] = 30'h1FE45982;
		ln_c_0[168] = 30'h1FD10763;
		ln_c_0[169] = 30'h1FBDC0E7;
		ln_c_0[170] = 30'h1FAA8600;
		ln_c_0[171] = 30'h1F9756A0;
		ln_c_0[172] = 30'h1F8432BB;
		ln_c_0[173] = 30'h1F711A42;
		ln_c_0[174] = 30'h1F5E0D26;
		ln_c_0[175] = 30'h1F4B0B5C;
		ln_c_0[176] = 30'h1F3814D4;
		ln_c_0[177] = 30'h1F252985;
		ln_c_0[178] = 30'h1F12495D;
		ln_c_0[179] = 30'h1EFF744E;
		ln_c_0[180] = 30'h1EECAA51;
		ln_c_0[181] = 30'h1ED9EB53;
		ln_c_0[182] = 30'h1EC7374D;
		ln_c_0[183] = 30'h1EB48E30;
		ln_c_0[184] = 30'h1EA1EFEB;
		ln_c_0[185] = 30'h1E8F5C76;
		ln_c_0[186] = 30'h1E7CD3C4;
		ln_c_0[187] = 30'h1E6A55C8;
		ln_c_0[188] = 30'h1E57E276;
		ln_c_0[189] = 30'h1E4579BF;
		ln_c_0[190] = 30'h1E331B9D;
		ln_c_0[191] = 30'h1E20C7FB;
		ln_c_0[192] = 30'h1E0E7ED5;
		ln_c_0[193] = 30'h1DFC401B;
		ln_c_0[194] = 30'h1DEA0BC2;
		ln_c_0[195] = 30'h1DD7E1BC;
		ln_c_0[196] = 30'h1DC5C203;
		ln_c_0[197] = 30'h1DB3AC88;
		ln_c_0[198] = 30'h1DA1A13F;
		ln_c_0[199] = 30'h1D8FA01C;
		ln_c_0[200] = 30'h1D7DA917;
		ln_c_0[201] = 30'h1D6BBC24;
		ln_c_0[202] = 30'h1D59D931;
		ln_c_0[203] = 30'h1D480038;
		ln_c_0[204] = 30'h1D36312F;
		ln_c_0[205] = 30'h1D246C0D;
		ln_c_0[206] = 30'h1D12B0BF;
		ln_c_0[207] = 30'h1D00FF41;
		ln_c_0[208] = 30'h1CEF5785;
		ln_c_0[209] = 30'h1CDDB981;
		ln_c_0[210] = 30'h1CCC252C;
		ln_c_0[211] = 30'h1CBA9A7A;
		ln_c_0[212] = 30'h1CA91960;
		ln_c_0[213] = 30'h1C97A1D7;
		ln_c_0[214] = 30'h1C8633CD;
		ln_c_0[215] = 30'h1C74CF3C;
		ln_c_0[216] = 30'h1C63741B;
		ln_c_0[217] = 30'h1C522260;
		ln_c_0[218] = 30'h1C40D9FF;
		ln_c_0[219] = 30'h1C2F9AED;
		ln_c_0[220] = 30'h1C1E6526;
		ln_c_0[221] = 30'h1C0D3897;
		ln_c_0[222] = 30'h1BFC153D;
		ln_c_0[223] = 30'h1BEAFB0A;
		ln_c_0[224] = 30'h1BD9E9F9;
		ln_c_0[225] = 30'h1BC8E1F9;
		ln_c_0[226] = 30'h1BB7E309;
		ln_c_0[227] = 30'h1BA6ED19;
		ln_c_0[228] = 30'h1B960023;
		ln_c_0[229] = 30'h1B851C1B;
		ln_c_0[230] = 30'h1B7440FB;
		ln_c_0[231] = 30'h1B636EB2;
		ln_c_0[232] = 30'h1B52A540;
		ln_c_0[233] = 30'h1B41E497;
		ln_c_0[234] = 30'h1B312CAB;
		ln_c_0[235] = 30'h1B207D7D;
		ln_c_0[236] = 30'h1B0FD6F8;
		ln_c_0[237] = 30'h1AFF391C;
		ln_c_0[238] = 30'h1AEEA3D8;
		ln_c_0[239] = 30'h1ADE172D;
		ln_c_0[240] = 30'h1ACD930B;
		ln_c_0[241] = 30'h1ABD176A;
		ln_c_0[242] = 30'h1AACA445;
		ln_c_0[243] = 30'h1A9C398C;
		ln_c_0[244] = 30'h1A8BD73D;
		ln_c_0[245] = 30'h1A7B7D4D;
		ln_c_0[246] = 30'h1A6B2BB3;
		ln_c_0[247] = 30'h1A5AE268;
		ln_c_0[248] = 30'h1A4AA167;
		ln_c_0[249] = 30'h1A3A689D;
		ln_c_0[250] = 30'h1A2A3803;
		ln_c_0[251] = 30'h1A1A0F9E;
		ln_c_0[252] = 30'h1A09EF5F;
		ln_c_0[253] = 30'h19F9D737;
		ln_c_0[254] = 30'h19E9C725;
		ln_c_0[255] = 30'h19D9BF23;
		
		c_0_t = ln_c_0[table_address_p1];
		c_1 = ln_c_1[table_address_p1];
		c_2 = ln_c_2[table_address_p1];
	end
//reset = 1? initialize all registers	
	if(reset != 1'b0)
	begin
		log_2_2 = 32'h0;
		value_d = 31'h0;
		expo_corr_d = 38'h0;
		leading_zeros_d = 6'h0;
		num2_d = 48'h0;
        temp_d = 30'h0;
        temp2_d = 30'h0;
		expo_d1 = 6'h0;
		expo_d2 = 6'h0;
		expo_d3 = 6'h0;
		expo_d4 = 6'h0;
		expo_d5 = 6'h0;
		expo_d6 = 6'h0;
		expo_d7 = 6'h0;
		mul2_d1 = 51'h0;
		mul2_d2 = 51'h0;
		mul3_d = 48'h0;
		mul3_t_d = 48'h0;
		t1_d = 30'h0;
		t2_d = 29'h0;
		t5_d = 28'h0;
		t1_d1 = 30'h0;
		t3_d1 = 30'h0;
		c_0_t_d1 = 19'h0;
		c_0_t_d2 = 19'h0;
		c_1_d1 = 22'h0;
		c_2_d1 = 30'h0;
		c_1_d2 = 22'h0;
        c_2_d2 = 30'h0;
		c_0_d1 = 19'h0;
		c_0_d2 = 19'h0;
		adj_log_val_d = 34'h0;
		shortened_num_d1 = 29'h0;
		shortened_num_d2 = 29'h0;
		shortened_num_d3 = 29'h0;
		shortened_num_d4 = 29'h0;
		shortened_num_dd1 = 29'h0;
		table_address_d1 = 8'h0;
		mul1_d = 29'h0;
		c_0_t = 19'h0;
		c_1 = 22'h0;
		c_2 = 30'h0;
		ln_c_2[0] = 19'h0;
		ln_c_2[1] = 19'h0;
		ln_c_2[2] = 19'h0;
		ln_c_2[3] = 19'h0;
		ln_c_2[4] = 19'h0;
		ln_c_2[5] = 19'h0;
		ln_c_2[6] = 19'h0;
		ln_c_2[7] = 19'h0;
		ln_c_2[8] = 19'h0;
		ln_c_2[9] = 19'h0;
		ln_c_2[10] = 19'h0;
		ln_c_2[11] = 19'h0;
		ln_c_2[12] = 19'h0;
		ln_c_2[13] = 19'h0;
		ln_c_2[14] = 19'h0;
		ln_c_2[15] = 19'h0;
		ln_c_2[16] = 19'h0;
		ln_c_2[17] = 19'h0;
		ln_c_2[18] = 19'h0;
		ln_c_2[19] = 19'h0;
		ln_c_2[20] = 19'h0;
		ln_c_2[21] = 19'h0;
		ln_c_2[22] = 19'h0;
		ln_c_2[23] = 19'h0;
		ln_c_2[24] = 19'h0;
		ln_c_2[25] = 19'h0;
		ln_c_2[26] = 19'h0;
		ln_c_2[27] = 19'h0;
		ln_c_2[28] = 19'h0;
		ln_c_2[29] = 19'h0;
		ln_c_2[30] = 19'h0;
		ln_c_2[31] = 19'h0;
		ln_c_2[32] = 19'h0;
		ln_c_2[33] = 19'h0;
		ln_c_2[34] = 19'h0;
		ln_c_2[35] = 19'h0;
		ln_c_2[36] = 19'h0;
		ln_c_2[37] = 19'h0;
		ln_c_2[38] = 19'h0;
		ln_c_2[39] = 19'h0;
		ln_c_2[40] = 19'h0;
		ln_c_2[41] = 19'h0;
		ln_c_2[42] = 19'h0;
		ln_c_2[43] = 19'h0;
		ln_c_2[44] = 19'h0;
		ln_c_2[45] = 19'h0;
		ln_c_2[46] = 19'h0;
		ln_c_2[47] = 19'h0;
		ln_c_2[48] = 19'h0;
		ln_c_2[49] = 19'h0;
		ln_c_2[50] = 19'h0;
		ln_c_2[51] = 19'h0;
		ln_c_2[52] = 19'h0;
		ln_c_2[53] = 19'h0;
		ln_c_2[54] = 19'h0;
		ln_c_2[55] = 19'h0;
		ln_c_2[56] = 19'h0;
		ln_c_2[57] = 19'h0;
		ln_c_2[58] = 19'h0;
		ln_c_2[59] = 19'h0;
		ln_c_2[60] = 19'h0;
		ln_c_2[61] = 19'h0;
		ln_c_2[62] = 19'h0;
		ln_c_2[63] = 19'h0;
		ln_c_2[64] = 19'h0;
		ln_c_2[65] = 19'h0;
		ln_c_2[66] = 19'h0;
		ln_c_2[67] = 19'h0;
		ln_c_2[68] = 19'h0;
		ln_c_2[69] = 19'h0;
		ln_c_2[70] = 19'h0;
		ln_c_2[71] = 19'h0;
		ln_c_2[72] = 19'h0;
		ln_c_2[73] = 19'h0;
		ln_c_2[74] = 19'h0;
		ln_c_2[75] = 19'h0;
		ln_c_2[76] = 19'h0;
		ln_c_2[77] = 19'h0;
		ln_c_2[78] = 19'h0;
		ln_c_2[79] = 19'h0;
		ln_c_2[80] = 19'h0;
		ln_c_2[81] = 19'h0;
		ln_c_2[82] = 19'h0;
		ln_c_2[83] = 19'h0;
		ln_c_2[84] = 19'h0;
		ln_c_2[85] = 19'h0;
		ln_c_2[86] = 19'h0;
		ln_c_2[87] = 19'h0;
		ln_c_2[88] = 19'h0;
		ln_c_2[89] = 19'h0;
		ln_c_2[90] = 19'h0;
		ln_c_2[91] = 19'h0;
		ln_c_2[92] = 19'h0;
		ln_c_2[93] = 19'h0;
		ln_c_2[94] = 19'h0;
		ln_c_2[95] = 19'h0;
		ln_c_2[96] = 19'h0;
		ln_c_2[97] = 19'h0;
		ln_c_2[98] = 19'h0;
		ln_c_2[99] = 19'h0;
		ln_c_2[100] = 19'h0;
		ln_c_2[101] = 19'h0;
		ln_c_2[102] = 19'h0;
		ln_c_2[103] = 19'h0;
		ln_c_2[104] = 19'h0;
		ln_c_2[105] = 19'h0;
		ln_c_2[106] = 19'h0;
		ln_c_2[107] = 19'h0;
		ln_c_2[108] = 19'h0;
		ln_c_2[109] = 19'h0;
		ln_c_2[110] = 19'h0;
		ln_c_2[111] = 19'h0;
		ln_c_2[112] = 19'h0;
		ln_c_2[113] = 19'h0;
		ln_c_2[114] = 19'h0;
		ln_c_2[115] = 19'h0;
		ln_c_2[116] = 19'h0;
		ln_c_2[117] = 19'h0;
		ln_c_2[118] = 19'h0;
		ln_c_2[119] = 19'h0;
		ln_c_2[120] = 19'h0;
		ln_c_2[121] = 19'h0;
		ln_c_2[122] = 19'h0;
		ln_c_2[123] = 19'h0;
		ln_c_2[124] = 19'h0;
		ln_c_2[125] = 19'h0;
		ln_c_2[126] = 19'h0;
		ln_c_2[127] = 19'h0;
		ln_c_2[128] = 19'h0;
		ln_c_2[129] = 19'h0;
		ln_c_2[130] = 19'h0;
		ln_c_2[131] = 19'h0;
		ln_c_2[132] = 19'h0;
		ln_c_2[133] = 19'h0;
		ln_c_2[134] = 19'h0;
		ln_c_2[135] = 19'h0;
		ln_c_2[136] = 19'h0;
		ln_c_2[137] = 19'h0;
		ln_c_2[138] = 19'h0;
		ln_c_2[139] = 19'h0;
		ln_c_2[140] = 19'h0;
		ln_c_2[141] = 19'h0;
		ln_c_2[142] = 19'h0;
		ln_c_2[143] = 19'h0;
		ln_c_2[144] = 19'h0;
		ln_c_2[145] = 19'h0;
		ln_c_2[146] = 19'h0;
		ln_c_2[147] = 19'h0;
		ln_c_2[148] = 19'h0;
		ln_c_2[149] = 19'h0;
		ln_c_2[150] = 19'h0;
		ln_c_2[151] = 19'h0;
		ln_c_2[152] = 19'h0;
		ln_c_2[153] = 19'h0;
		ln_c_2[154] = 19'h0;
		ln_c_2[155] = 19'h0;
		ln_c_2[156] = 19'h0;
		ln_c_2[157] = 19'h0;
		ln_c_2[158] = 19'h0;
		ln_c_2[159] = 19'h0;
		ln_c_2[160] = 19'h0;
		ln_c_2[161] = 19'h0;
		ln_c_2[162] = 19'h0;
		ln_c_2[163] = 19'h0;
		ln_c_2[164] = 19'h0;
		ln_c_2[165] = 19'h0;
		ln_c_2[166] = 19'h0;
		ln_c_2[167] = 19'h0;
		ln_c_2[168] = 19'h0;
		ln_c_2[169] = 19'h0;
		ln_c_2[170] = 19'h0;
		ln_c_2[171] = 19'h0;
		ln_c_2[172] = 19'h0;
		ln_c_2[173] = 19'h0;
		ln_c_2[174] = 19'h0;
		ln_c_2[175] = 19'h0;
		ln_c_2[176] = 19'h0;
		ln_c_2[177] = 19'h0;
		ln_c_2[178] = 19'h0;
		ln_c_2[179] = 19'h0;
		ln_c_2[180] = 19'h0;
		ln_c_2[181] = 19'h0;
		ln_c_2[182] = 19'h0;
		ln_c_2[183] = 19'h0;
		ln_c_2[184] = 19'h0;
		ln_c_2[185] = 19'h0;
		ln_c_2[186] = 19'h0;
		ln_c_2[187] = 19'h0;
		ln_c_2[188] = 19'h0;
		ln_c_2[189] = 19'h0;
		ln_c_2[190] = 19'h0;
		ln_c_2[191] = 19'h0;
		ln_c_2[192] = 19'h0;
		ln_c_2[193] = 19'h0;
		ln_c_2[194] = 19'h0;
		ln_c_2[195] = 19'h0;
		ln_c_2[196] = 19'h0;
		ln_c_2[197] = 19'h0;
		ln_c_2[198] = 19'h0;
		ln_c_2[199] = 19'h0;
		ln_c_2[200] = 19'h0;
		ln_c_2[201] = 19'h0;
		ln_c_2[202] = 19'h0;
		ln_c_2[203] = 19'h0;
		ln_c_2[204] = 19'h0;
		ln_c_2[205] = 19'h0;
		ln_c_2[206] = 19'h0;
		ln_c_2[207] = 19'h0;
		ln_c_2[208] = 19'h0;
		ln_c_2[209] = 19'h0;
		ln_c_2[210] = 19'h0;
		ln_c_2[211] = 19'h0;
		ln_c_2[212] = 19'h0;
		ln_c_2[213] = 19'h0;
		ln_c_2[214] = 19'h0;
		ln_c_2[215] = 19'h0;
		ln_c_2[216] = 19'h0;
		ln_c_2[217] = 19'h0;
		ln_c_2[218] = 19'h0;
		ln_c_2[219] = 19'h0;
		ln_c_2[220] = 19'h0;
		ln_c_2[221] = 19'h0;
		ln_c_2[222] = 19'h0;
		ln_c_2[223] = 19'h0;
		ln_c_2[224] = 19'h0;
		ln_c_2[225] = 19'h0;
		ln_c_2[226] = 19'h0;
		ln_c_2[227] = 19'h0;
		ln_c_2[228] = 19'h0;
		ln_c_2[229] = 19'h0;
		ln_c_2[230] = 19'h0;
		ln_c_2[231] = 19'h0;
		ln_c_2[232] = 19'h0;
		ln_c_2[233] = 19'h0;
		ln_c_2[234] = 19'h0;
		ln_c_2[235] = 19'h0;
		ln_c_2[236] = 19'h0;
		ln_c_2[237] = 19'h0;
		ln_c_2[238] = 19'h0;
		ln_c_2[239] = 19'h0;
		ln_c_2[240] = 19'h0;
		ln_c_2[241] = 19'h0;
		ln_c_2[242] = 19'h0;
		ln_c_2[243] = 19'h0;
		ln_c_2[244] = 19'h0;
		ln_c_2[245] = 19'h0;
		ln_c_2[246] = 19'h0;
		ln_c_2[247] = 19'h0;
		ln_c_2[248] = 19'h0;
		ln_c_2[249] = 19'h0;
		ln_c_2[250] = 19'h0;
		ln_c_2[251] = 19'h0;
		ln_c_2[252] = 19'h0;
		ln_c_2[253] = 19'h0;
		ln_c_2[254] = 19'h0;
		ln_c_2[255] = 19'h0;

		ln_c_1[0] = 22'h0;
		ln_c_1[1] = 22'h0;
		ln_c_1[2] = 22'h0;
		ln_c_1[3] = 22'h0;
		ln_c_1[4] = 22'h0;
		ln_c_1[5] = 22'h0;
		ln_c_1[6] = 22'h0;
		ln_c_1[7] = 22'h0;
		ln_c_1[8] = 22'h0;
		ln_c_1[9] = 22'h0;
		ln_c_1[10] = 22'h0;
		ln_c_1[11] = 22'h0;
		ln_c_1[12] = 22'h0;
		ln_c_1[13] = 22'h0;
		ln_c_1[14] = 22'h0;
		ln_c_1[15] = 22'h0;
		ln_c_1[16] = 22'h0;
		ln_c_1[17] = 22'h0;
		ln_c_1[18] = 22'h0;
		ln_c_1[19] = 22'h0;
		ln_c_1[20] = 22'h0;
		ln_c_1[21] = 22'h0;
		ln_c_1[22] = 22'h0;
		ln_c_1[23] = 22'h0;
		ln_c_1[24] = 22'h0;
		ln_c_1[25] = 22'h0;
		ln_c_1[26] = 22'h0;
		ln_c_1[27] = 22'h0;
		ln_c_1[28] = 22'h0;
		ln_c_1[29] = 22'h0;
		ln_c_1[30] = 22'h0;
		ln_c_1[31] = 22'h0;
		ln_c_1[32] = 22'h0;
		ln_c_1[33] = 22'h0;
		ln_c_1[34] = 22'h0;
		ln_c_1[35] = 22'h0;
		ln_c_1[36] = 22'h0;
		ln_c_1[37] = 22'h0;
		ln_c_1[38] = 22'h0;
		ln_c_1[39] = 22'h0;
		ln_c_1[40] = 22'h0;
		ln_c_1[41] = 22'h0;
		ln_c_1[42] = 22'h0;
		ln_c_1[43] = 22'h0;
		ln_c_1[44] = 22'h0;
		ln_c_1[45] = 22'h0;
		ln_c_1[46] = 22'h0;
		ln_c_1[47] = 22'h0;
		ln_c_1[48] = 22'h0;
		ln_c_1[49] = 22'h0;
		ln_c_1[50] = 22'h0;
		ln_c_1[51] = 22'h0;
		ln_c_1[52] = 22'h0;
		ln_c_1[53] = 22'h0;
		ln_c_1[54] = 22'h0;
		ln_c_1[55] = 22'h0;
		ln_c_1[56] = 22'h0;
		ln_c_1[57] = 22'h0;
		ln_c_1[58] = 22'h0;
		ln_c_1[59] = 22'h0;
		ln_c_1[60] = 22'h0;
		ln_c_1[61] = 22'h0;
		ln_c_1[62] = 22'h0;
		ln_c_1[63] = 22'h0;
		ln_c_1[64] = 22'h0;
		ln_c_1[65] = 22'h0;
		ln_c_1[66] = 22'h0;
		ln_c_1[67] = 22'h0;
		ln_c_1[68] = 22'h0;
		ln_c_1[69] = 22'h0;
		ln_c_1[70] = 22'h0;
		ln_c_1[71] = 22'h0;
		ln_c_1[72] = 22'h0;
		ln_c_1[73] = 22'h0;
		ln_c_1[74] = 22'h0;
		ln_c_1[75] = 22'h0;
		ln_c_1[76] = 22'h0;
		ln_c_1[77] = 22'h0;
		ln_c_1[78] = 22'h0;
		ln_c_1[79] = 22'h0;
		ln_c_1[80] = 22'h0;
		ln_c_1[81] = 22'h0;
		ln_c_1[82] = 22'h0;
		ln_c_1[83] = 22'h0;
		ln_c_1[84] = 22'h0;
		ln_c_1[85] = 22'h0;
		ln_c_1[86] = 22'h0;
		ln_c_1[87] = 22'h0;
		ln_c_1[88] = 22'h0;
		ln_c_1[89] = 22'h0;
		ln_c_1[90] = 22'h0;
		ln_c_1[91] = 22'h0;
		ln_c_1[92] = 22'h0;
		ln_c_1[93] = 22'h0;
		ln_c_1[94] = 22'h0;
		ln_c_1[95] = 22'h0;
		ln_c_1[96] = 22'h0;
		ln_c_1[97] = 22'h0;
		ln_c_1[98] = 22'h0;
		ln_c_1[99] = 22'h0;
		ln_c_1[100] = 22'h0;
		ln_c_1[101] = 22'h0;
		ln_c_1[102] = 22'h0;
		ln_c_1[103] = 22'h0;
		ln_c_1[104] = 22'h0;
		ln_c_1[105] = 22'h0;
		ln_c_1[106] = 22'h0;
		ln_c_1[107] = 22'h0;
		ln_c_1[108] = 22'h0;
		ln_c_1[109] = 22'h0;
		ln_c_1[110] = 22'h0;
		ln_c_1[111] = 22'h0;
		ln_c_1[112] = 22'h0;
		ln_c_1[113] = 22'h0;
		ln_c_1[114] = 22'h0;
		ln_c_1[115] = 22'h0;
		ln_c_1[116] = 22'h0;
		ln_c_1[117] = 22'h0;
		ln_c_1[118] = 22'h0;
		ln_c_1[119] = 22'h0;
		ln_c_1[120] = 22'h0;
		ln_c_1[121] = 22'h0;
		ln_c_1[122] = 22'h0;
		ln_c_1[123] = 22'h0;
		ln_c_1[124] = 22'h0;
		ln_c_1[125] = 22'h0;
		ln_c_1[126] = 22'h0;
		ln_c_1[127] = 22'h0;
		ln_c_1[128] = 22'h0;
		ln_c_1[129] = 22'h0;
		ln_c_1[130] = 22'h0;
		ln_c_1[131] = 22'h0;
		ln_c_1[132] = 22'h0;
		ln_c_1[133] = 22'h0;
		ln_c_1[134] = 22'h0;
		ln_c_1[135] = 22'h0;
		ln_c_1[136] = 22'h0;
		ln_c_1[137] = 22'h0;
		ln_c_1[138] = 22'h0;
		ln_c_1[139] = 22'h0;
		ln_c_1[140] = 22'h0;
		ln_c_1[141] = 22'h0;
		ln_c_1[142] = 22'h0;
		ln_c_1[143] = 22'h0;
		ln_c_1[144] = 22'h0;
		ln_c_1[145] = 22'h0;
		ln_c_1[146] = 22'h0;
		ln_c_1[147] = 22'h0;
		ln_c_1[148] = 22'h0;
		ln_c_1[149] = 22'h0;
		ln_c_1[150] = 22'h0;
		ln_c_1[151] = 22'h0;
		ln_c_1[152] = 22'h0;
		ln_c_1[153] = 22'h0;
		ln_c_1[154] = 22'h0;
		ln_c_1[155] = 22'h0;
		ln_c_1[156] = 22'h0;
		ln_c_1[157] = 22'h0;
		ln_c_1[158] = 22'h0;
		ln_c_1[159] = 22'h0;
		ln_c_1[160] = 22'h0;
		ln_c_1[161] = 22'h0;
		ln_c_1[162] = 22'h0;
		ln_c_1[163] = 22'h0;
		ln_c_1[164] = 22'h0;
		ln_c_1[165] = 22'h0;
		ln_c_1[166] = 22'h0;
		ln_c_1[167] = 22'h0;
		ln_c_1[168] = 22'h0;
		ln_c_1[169] = 22'h0;
		ln_c_1[170] = 22'h0;
		ln_c_1[171] = 22'h0;
		ln_c_1[172] = 22'h0;
		ln_c_1[173] = 22'h0;
		ln_c_1[174] = 22'h0;
		ln_c_1[175] = 22'h0;
		ln_c_1[176] = 22'h0;
		ln_c_1[177] = 22'h0;
		ln_c_1[178] = 22'h0;
		ln_c_1[179] = 22'h0;
		ln_c_1[180] = 22'h0;
		ln_c_1[181] = 22'h0;
		ln_c_1[182] = 22'h0;
		ln_c_1[183] = 22'h0;
		ln_c_1[184] = 22'h0;
		ln_c_1[185] = 22'h0;
		ln_c_1[186] = 22'h0;
		ln_c_1[187] = 22'h0;
		ln_c_1[188] = 22'h0;
		ln_c_1[189] = 22'h0;
		ln_c_1[190] = 22'h0;
		ln_c_1[191] = 22'h0;
		ln_c_1[192] = 22'h0;
		ln_c_1[193] = 22'h0;
		ln_c_1[194] = 22'h0;
		ln_c_1[195] = 22'h0;
		ln_c_1[196] = 22'h0;
		ln_c_1[197] = 22'h0;
		ln_c_1[198] = 22'h0;
		ln_c_1[199] = 22'h0;
		ln_c_1[200] = 22'h0;
		ln_c_1[201] = 22'h0;
		ln_c_1[202] = 22'h0;
		ln_c_1[203] = 22'h0;
		ln_c_1[204] = 22'h0;
		ln_c_1[205] = 22'h0;
		ln_c_1[206] = 22'h0;
		ln_c_1[207] = 22'h0;
		ln_c_1[208] = 22'h0;
		ln_c_1[209] = 22'h0;
		ln_c_1[210] = 22'h0;
		ln_c_1[211] = 22'h0;
		ln_c_1[212] = 22'h0;
		ln_c_1[213] = 22'h0;
		ln_c_1[214] = 22'h0;
		ln_c_1[215] = 22'h0;
		ln_c_1[216] = 22'h0;
		ln_c_1[217] = 22'h0;
		ln_c_1[218] = 22'h0;
		ln_c_1[219] = 22'h0;
		ln_c_1[220] = 22'h0;
		ln_c_1[221] = 22'h0;
		ln_c_1[222] = 22'h0;
		ln_c_1[223] = 22'h0;
		ln_c_1[224] = 22'h0;
		ln_c_1[225] = 22'h0;
		ln_c_1[226] = 22'h0;
		ln_c_1[227] = 22'h0;
		ln_c_1[228] = 22'h0;
		ln_c_1[229] = 22'h0;
		ln_c_1[230] = 22'h0;
		ln_c_1[231] = 22'h0;
		ln_c_1[232] = 22'h0;
		ln_c_1[233] = 22'h0;
		ln_c_1[234] = 22'h0;
		ln_c_1[235] = 22'h0;
		ln_c_1[236] = 22'h0;
		ln_c_1[237] = 22'h0;
		ln_c_1[238] = 22'h0;
		ln_c_1[239] = 22'h0;
		ln_c_1[240] = 22'h0;
		ln_c_1[241] = 22'h0;
		ln_c_1[242] = 22'h0;
		ln_c_1[243] = 22'h0;
		ln_c_1[244] = 22'h0;
		ln_c_1[245] = 22'h0;
		ln_c_1[246] = 22'h0;
		ln_c_1[247] = 22'h0;
		ln_c_1[248] = 22'h0;
		ln_c_1[249] = 22'h0;
		ln_c_1[250] = 22'h0;
		ln_c_1[251] = 22'h0;
		ln_c_1[252] = 22'h0;
		ln_c_1[253] = 22'h0;
		ln_c_1[254] = 22'h0;
		ln_c_1[255] = 22'h0;

		ln_c_0[0] = 30'h0;
		ln_c_0[1] = 30'h0;
		ln_c_0[2] = 30'h0;
		ln_c_0[3] = 30'h0;
		ln_c_0[4] = 30'h0;
		ln_c_0[5] = 30'h0;
		ln_c_0[6] = 30'h0;
		ln_c_0[7] = 30'h0;
		ln_c_0[8] = 30'h0;
		ln_c_0[9] = 30'h0;
		ln_c_0[10] = 30'h0;
		ln_c_0[11] = 30'h0;
		ln_c_0[12] = 30'h0;
		ln_c_0[13] = 30'h0;
		ln_c_0[14] = 30'h0;
		ln_c_0[15] = 30'h0;
		ln_c_0[16] = 30'h0;
		ln_c_0[17] = 30'h0;
		ln_c_0[18] = 30'h0;
		ln_c_0[19] = 30'h0;
		ln_c_0[20] = 30'h0;
		ln_c_0[21] = 30'h0;
		ln_c_0[22] = 30'h0;
		ln_c_0[23] = 30'h0;
		ln_c_0[24] = 30'h0;
		ln_c_0[25] = 30'h0;
		ln_c_0[26] = 30'h0;
		ln_c_0[27] = 30'h0;
		ln_c_0[28] = 30'h0;
		ln_c_0[29] = 30'h0;
		ln_c_0[30] = 30'h0;
		ln_c_0[31] = 30'h0;
		ln_c_0[32] = 30'h0;
		ln_c_0[33] = 30'h0;
		ln_c_0[34] = 30'h0;
		ln_c_0[35] = 30'h0;
		ln_c_0[36] = 30'h0;
		ln_c_0[37] = 30'h0;
		ln_c_0[38] = 30'h0;
		ln_c_0[39] = 30'h0;
		ln_c_0[40] = 30'h0;
		ln_c_0[41] = 30'h0;
		ln_c_0[42] = 30'h0;
		ln_c_0[43] = 30'h0;
		ln_c_0[44] = 30'h0;
		ln_c_0[45] = 30'h0;
		ln_c_0[46] = 30'h0;
		ln_c_0[47] = 30'h0;
		ln_c_0[48] = 30'h0;
		ln_c_0[49] = 30'h0;
		ln_c_0[50] = 30'h0;
		ln_c_0[51] = 30'h0;
		ln_c_0[52] = 30'h0;
		ln_c_0[53] = 30'h0;
		ln_c_0[54] = 30'h0;
		ln_c_0[55] = 30'h0;
		ln_c_0[56] = 30'h0;
		ln_c_0[57] = 30'h0;
		ln_c_0[58] = 30'h0;
		ln_c_0[59] = 30'h0;
		ln_c_0[60] = 30'h0;
		ln_c_0[61] = 30'h0;
		ln_c_0[62] = 30'h0;
		ln_c_0[63] = 30'h0;
		ln_c_0[64] = 30'h0;
		ln_c_0[65] = 30'h0;
		ln_c_0[66] = 30'h0;
		ln_c_0[67] = 30'h0;
		ln_c_0[68] = 30'h0;
		ln_c_0[69] = 30'h0;
		ln_c_0[70] = 30'h0;
		ln_c_0[71] = 30'h0;
		ln_c_0[72] = 30'h0;
		ln_c_0[73] = 30'h0;
		ln_c_0[74] = 30'h0;
		ln_c_0[75] = 30'h0;
		ln_c_0[76] = 30'h0;
		ln_c_0[77] = 30'h0;
		ln_c_0[78] = 30'h0;
		ln_c_0[79] = 30'h0;
		ln_c_0[80] = 30'h0;
		ln_c_0[81] = 30'h0;
		ln_c_0[82] = 30'h0;
		ln_c_0[83] = 30'h0;
		ln_c_0[84] = 30'h0;
		ln_c_0[85] = 30'h0;
		ln_c_0[86] = 30'h0;
		ln_c_0[87] = 30'h0;
		ln_c_0[88] = 30'h0;
		ln_c_0[89] = 30'h0;
		ln_c_0[90] = 30'h0;
		ln_c_0[91] = 30'h0;
		ln_c_0[92] = 30'h0;
		ln_c_0[93] = 30'h0;
		ln_c_0[94] = 30'h0;
		ln_c_0[95] = 30'h0;
		ln_c_0[96] = 30'h0;
		ln_c_0[97] = 30'h0;
		ln_c_0[98] = 30'h0;
		ln_c_0[99] = 30'h0;
		ln_c_0[100] = 30'h0;
		ln_c_0[101] = 30'h0;
		ln_c_0[102] = 30'h0;
		ln_c_0[103] = 30'h0;
		ln_c_0[104] = 30'h0;
		ln_c_0[105] = 30'h0;
		ln_c_0[106] = 30'h0;
		ln_c_0[107] = 30'h0;
		ln_c_0[108] = 30'h0;
		ln_c_0[109] = 30'h0;
		ln_c_0[110] = 30'h0;
		ln_c_0[111] = 30'h0;
		ln_c_0[112] = 30'h0;
		ln_c_0[113] = 30'h0;
		ln_c_0[114] = 30'h0;
		ln_c_0[115] = 30'h0;
		ln_c_0[116] = 30'h0;
		ln_c_0[117] = 30'h0;
		ln_c_0[118] = 30'h0;
		ln_c_0[119] = 30'h0;
		ln_c_0[120] = 30'h0;
		ln_c_0[121] = 30'h0;
		ln_c_0[122] = 30'h0;
		ln_c_0[123] = 30'h0;
		ln_c_0[124] = 30'h0;
		ln_c_0[125] = 30'h0;
		ln_c_0[126] = 30'h0;
		ln_c_0[127] = 30'h0;
		ln_c_0[128] = 30'h0;
		ln_c_0[129] = 30'h0;
		ln_c_0[130] = 30'h0;
		ln_c_0[131] = 30'h0;
		ln_c_0[132] = 30'h0;
		ln_c_0[133] = 30'h0;
		ln_c_0[134] = 30'h0;
		ln_c_0[135] = 30'h0;
		ln_c_0[136] = 30'h0;
		ln_c_0[137] = 30'h0;
		ln_c_0[138] = 30'h0;
		ln_c_0[139] = 30'h0;
		ln_c_0[140] = 30'h0;
		ln_c_0[141] = 30'h0;
		ln_c_0[142] = 30'h0;
		ln_c_0[143] = 30'h0;
		ln_c_0[144] = 30'h0;
		ln_c_0[145] = 30'h0;
		ln_c_0[146] = 30'h0;
		ln_c_0[147] = 30'h0;
		ln_c_0[148] = 30'h0;
		ln_c_0[149] = 30'h0;
		ln_c_0[150] = 30'h0;
		ln_c_0[151] = 30'h0;
		ln_c_0[152] = 30'h0;
		ln_c_0[153] = 30'h0;
		ln_c_0[154] = 30'h0;
		ln_c_0[155] = 30'h0;
		ln_c_0[156] = 30'h0;
		ln_c_0[157] = 30'h0;
		ln_c_0[158] = 30'h0;
		ln_c_0[159] = 30'h0;
		ln_c_0[160] = 30'h0;
		ln_c_0[161] = 30'h0;
		ln_c_0[162] = 30'h0;
		ln_c_0[163] = 30'h0;
		ln_c_0[164] = 30'h0;
		ln_c_0[165] = 30'h0;
		ln_c_0[166] = 30'h0;
		ln_c_0[167] = 30'h0;
		ln_c_0[168] = 30'h0;
		ln_c_0[169] = 30'h0;
		ln_c_0[170] = 30'h0;
		ln_c_0[171] = 30'h0;
		ln_c_0[172] = 30'h0;
		ln_c_0[173] = 30'h0;
		ln_c_0[174] = 30'h0;
		ln_c_0[175] = 30'h0;
		ln_c_0[176] = 30'h0;
		ln_c_0[177] = 30'h0;
		ln_c_0[178] = 30'h0;
		ln_c_0[179] = 30'h0;
		ln_c_0[180] = 30'h0;
		ln_c_0[181] = 30'h0;
		ln_c_0[182] = 30'h0;
		ln_c_0[183] = 30'h0;
		ln_c_0[184] = 30'h0;
		ln_c_0[185] = 30'h0;
		ln_c_0[186] = 30'h0;
		ln_c_0[187] = 30'h0;
		ln_c_0[188] = 30'h0;
		ln_c_0[189] = 30'h0;
		ln_c_0[190] = 30'h0;
		ln_c_0[191] = 30'h0;
		ln_c_0[192] = 30'h0;
		ln_c_0[193] = 30'h0;
		ln_c_0[194] = 30'h0;
		ln_c_0[195] = 30'h0;
		ln_c_0[196] = 30'h0;
		ln_c_0[197] = 30'h0;
		ln_c_0[198] = 30'h0;
		ln_c_0[199] = 30'h0;
		ln_c_0[200] = 30'h0;
		ln_c_0[201] = 30'h0;
		ln_c_0[202] = 30'h0;
		ln_c_0[203] = 30'h0;
		ln_c_0[204] = 30'h0;
		ln_c_0[205] = 30'h0;
		ln_c_0[206] = 30'h0;
		ln_c_0[207] = 30'h0;
		ln_c_0[208] = 30'h0;
		ln_c_0[209] = 30'h0;
		ln_c_0[210] = 30'h0;
		ln_c_0[211] = 30'h0;
		ln_c_0[212] = 30'h0;
		ln_c_0[213] = 30'h0;
		ln_c_0[214] = 30'h0;
		ln_c_0[215] = 30'h0;
		ln_c_0[216] = 30'h0;
		ln_c_0[217] = 30'h0;
		ln_c_0[218] = 30'h0;
		ln_c_0[219] = 30'h0;
		ln_c_0[220] = 30'h0;
		ln_c_0[221] = 30'h0;
		ln_c_0[222] = 30'h0;
		ln_c_0[223] = 30'h0;
		ln_c_0[224] = 30'h0;
		ln_c_0[225] = 30'h0;
		ln_c_0[226] = 30'h0;
		ln_c_0[227] = 30'h0;
		ln_c_0[228] = 30'h0;
		ln_c_0[229] = 30'h0;
		ln_c_0[230] = 30'h0;
		ln_c_0[231] = 30'h0;
		ln_c_0[232] = 30'h0;
		ln_c_0[233] = 30'h0;
		ln_c_0[234] = 30'h0;
		ln_c_0[235] = 30'h0;
		ln_c_0[236] = 30'h0;
		ln_c_0[237] = 30'h0;
		ln_c_0[238] = 30'h0;
		ln_c_0[239] = 30'h0;
		ln_c_0[240] = 30'h0;
		ln_c_0[241] = 30'h0;
		ln_c_0[242] = 30'h0;
		ln_c_0[243] = 30'h0;
		ln_c_0[244] = 30'h0;
		ln_c_0[245] = 30'h0;
		ln_c_0[246] = 30'h0;
		ln_c_0[247] = 30'h0;
		ln_c_0[248] = 30'h0;
		ln_c_0[249] = 30'h0;
		ln_c_0[250] = 30'h0;
		ln_c_0[251] = 30'h0;
		ln_c_0[252] = 30'h0;
		ln_c_0[253] = 30'h0;
		ln_c_0[254] = 30'h0;
		ln_c_0[255] = 30'h0;
	end
end

//end
endmodule